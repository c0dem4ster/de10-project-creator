-- name:    [project].vhd
-- author:  [author]
-- date:    [date]
-- content: [description]

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.math_real.all;

entity [project] is
  port(RESET_n : in std_logic;
       CLK     : in std_logic);
end [project];

architecture rtl of [project] is
begin
end rtl;